`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ece274a
// Engineer: Ali Akoglu 
// 
// Create Date:    21:12:26 04/09/2015 
// Design Name: 
// Module Name:    sort_TB 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sort_TB(    );

//DataMemory memory(t_d_add, t_wd_val, t_clk, t_s_dmw, t_s_dmr, t_rdata); 
reg Clk;
reg Go, Rst;

wire [4:0] Address;
wire [7:0] ReadData,WriteData;
wire MemRead,MemWrite;

integer i;

sort_top my_sort(Go, Rst, Clk, 8'd32, ReadData, Address, WriteData, MemWrite, MemRead);
DataMemory my_memory(Address, WriteData, Clk, MemWrite, MemRead, ReadData); 

/*
 Go, Rst, Clk, 32:  are the inputs to the sort top module generated by the testbench.
 						 here 32 is the array size. we will be sorting 32 elements
 ReadData: 
				8-bit data read from the memory
 Address: 
				datapath generates the 5-bit address to read from or write into the memory  
 WriteData: 
				datapath generates the 8-bit value to be written into the memory
 MemWrite, MemRead: 
				State machine enables the reads from the memory or writes into the memory and generates 
*/

// sort_top is the top module that integrates datapath and controller 
// use this exact name and port names and order 
// your top module receives 32 as an input. Make sure that your datapath works for any array size

always begin
	Clk <=1;
	#5;
	Clk<=0;
	#5;
end

initial begin
Rst <=1;
Go<=0;

@(posedge Clk);
#5;
Rst <=0;
Go <= 1;

@(posedge Clk);
#5;
Go <=0;

for (i=0; i<2000;i=i+1) begin
	@(posedge Clk);
	//#5;
	//Address <= i;
  
end
end
endmodule
